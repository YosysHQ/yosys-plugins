entity e1 is
    Port (
        a: in  STD_LOGIC;
        b,c,d: out  STD_LOGIC;
        e,f: in  STD_LOGIC
    );
end e1;
