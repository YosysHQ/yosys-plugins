entity e1 is
    Port (
        a: in  STD_LOGIC;
        b: out  STD_LOGIC
    );
end e1;
